module a;
x
endmodule
